\m5_TLV_version 1d: tl-x.org
\m5
   
   // ============================================
   // Welcome, new visitors! Try the "Learn" menu.
   // ============================================
   
   //use(m5-1.0)   /// uncomment to use M5 macro library.
\SV
   // Macro providing required top-level module definition, random
   // stimulus support, and Verilator config.
   m5_makerchip_module   // (Expanded in Nav-TLV pane.)
   //module andg(input in1,output out1);
   //out1 = in1;
   //endmodule

\TLV
   //$reset = *reset;
   
   //$out = ($sel==1'b0) ? $a : $b; 
   $out = $sel[1] ? ($sel[0] ? $d : $c) : ($sel[0] ? $b : $a) ; 
   
   // Assert these to end simulation (before the cycle limit).
   *passed = *cyc_cnt > 40;
   *failed = 1'b0;
\SV
   endmodule
